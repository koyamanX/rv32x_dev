../SDRAM_Controler/simulation/sdr_parameters.vh